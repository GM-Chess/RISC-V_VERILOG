module yAdder1(z, cout, a, b, cin);

    output z, cout;
    input a, b, cin;
    wire tmp, outR, outL;

    xor left_xor(tmp, a, b);
    xor right_xor(z, cin, tmp);
    and left_and(outL, cin, tmp);
    and right_and(outR, a, b);
    or anOR(cout, outL, outR);

endmodule 